`timescale 1ns/1ps

module Game_FSM(
	input                CLK,
	input                RESET,
	input      [2:0]     KEY_VALUE,
	input                KEY_VALID,
	output reg [4*9-1:0] CONTROL_ARRAY
);


endmodule